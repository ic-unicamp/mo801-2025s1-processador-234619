module clocked_register(
    input
)